D:\Nute\Armlet\Simulation\Twin-T Single-Op Band-Pass.CIR Transient,AC Analysis
* Spectrum Software Micro-Cap 9.0.7
* Date 27.10.2012 Time 18:07:27
* Converted From Micro Cap Source file to PSPICE
*
.FUNC DPWR(D) {I(D)*V(D)}
.FUNC BPWR(Q) {IC(Q)*VCE(Q)+IB(Q)*VBE(Q)}
.FUNC FPWR(M) {ID(M)*VDS(M)}
.FUNC HOTD(D,MAX) {IF((V(D)*I(D)>MAX),1,0)}
.FUNC HOTB(Q,MAX) {IF((VCE(Q)*IC(Q)+IB(Q)*VBE(Q)>MAX),1,0)}
.FUNC HOTF(M,MAX) {IF((VDS(M)*ID(M)>MAX),1,0)}
.PARAM LOW3MIN={IMPORT(LOW3MIN.OUT,LOW3THRES)}
.PARAM HIGH3MAX={IMPORT(HIGH3MAX.OUT,HIGH3THRES)}
.PARAM LOWLVDS={IMPORT(LOWLVDS.OUT,LOWLIMIT)}
.PARAM HILVDS={IMPORT(HILVDS.OUT,HILIMIT)}
.PARAM LIMTLVDS={IMPORT(LIMTLVDS.OUT,LVDSLIMITS)}
.FUNC SKINAC(DCRES,RESISTIVITY,RELPERM,RADIUS) {((PI*RADIUS*RADIUS)/((PI*RADIUS*RADIUS)-PI*(RADIUS-SKINDEPTHAC(RESISTIVITY,RELPERM))**2))*DCRES}
.FUNC SKINDEPTHAC(RESISTIVITY,RELPERM) {503.3*(SQRT(RESISTIVITY/(RELPERM*F)))}
.FUNC SKINTR(DCRES,RESISTIVITY,RELPERM,RADIUS,FREQ) {((PI*RADIUS*RADIUS)/((PI*RADIUS*RADIUS)-PI*(RADIUS-SKINDEPTHTR(RESISTIVITY,RELPERM,FREQ))**2))*DCRES}
.FUNC SKINDEPTHTR(RESISTIVITY,RELPERM,FREQ) {503.3*(SQRT(RESISTIVITY/(RELPERM*FREQ)))}
.PARAM FREQVAL=307KHZ
.PARAM RGAIN=10K
.PARAM CVAL=1000PF
.PARAM RVAL=1.5K
C1 5 7 {Cval}
C2 7 Out1 {Cval}
C3 6 Vcc/2 {Cval*2}
CIN Input 4 10u
CSH 3 0 0.1u
R1 5 6 {Rval}
R2 Out1 6 {Rval}
R3 7 Vcc/2 {Rval/2}
R4 10 4 {Rgain}
R5 Vcc/2 10 1k
RDOWN 0 3 100k
RUP 3 Vcc 100k
V1 INTERIOR_NONE1 0 AC 1 SIN (0 10MV FREQVAL 0 0 0)
RV1 Input INTERIOR_NONE1 2.5 ;added by V1
V2 Vcc 0 3.3V
X3 3 Vcc/2 Vcc 0 Vcc/2 AD8515
X4 10 5 Vcc 0 Out1 MC33174_MC
*
.OPTIONS ACCT LIST OPTS ABSTOL=1pA CHGTOL=.01pC DEFL=100u DEFW=100u DEFNRD=0
+ DEFNRS=0 DEFPD=0 DEFPS=0 DIGDRVF=2 DIGDRVZ=20K DIGERRDEFAULT=20 DIGERRLIMIT=0
+ DIGFREQ=10GHz DIGINITSTATE=0 DIGIOLVL=2 DIGMNTYMX=2 DIGMNTYSCALE=0.4 DIGOVRDRV=3
+ DIGTYMXSCALE=1.6 GMIN=1p ITL1=100 ITL2=50 ITL4=10 PIVREL=1m PIVTOL=.1p RELTOL=1m
+ TNOM=27 TRTOL=7 VNTOL=1u WIDTH=80
*
.LIB "C:\MC9\library\NOM.LIB"
*
.TEMP 27
*
.TRAN 3e-005 1.5m 0 
.PRINT TRAN V([INPUT])
.PLOT TRAN V([INPUT])
.PRINT TRAN V([OUT1])
.PLOT TRAN V([OUT1])
*
.AC LIN 29999 10kHz 300kHz
.PRINT AC VDB([OUT1])
.PLOT AC VDB([OUT1])
*
.PROBE
.END
;$SpiceType=PSPICE
